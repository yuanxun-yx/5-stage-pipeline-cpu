`ifndef DEBUG_VH
`define DEBUG_VH

//`define DEBUG_MODE

`endif